Common Emmitter o/p characteristics

Vcc 5 0 10V
Vbb 3 0 3V
Rc 2 5 2k
Rb 1 3 220k
Q1 2 1 0 Q2N2222

.dc Vbb 0 3 0.1V Vcc 10 0 2V 
.lib nom.lib
.probe 
.end

