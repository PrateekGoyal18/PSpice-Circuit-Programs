*FULL WAVE
 D1 0 1 D1N4002
D2 1 3 D1N4002
D3 2 3 D1N4002
D4 0 2 D1N4002
R1 0 3 1K

V1 1 2 SIN(1 10 100)

.TRAN 0.1m 50m 30m 0.1m
.PROBE
.END
