MOSFET characteristics Id v/s Vds

Vgs 1 0 4V
Vds 2 0 10V
M1 2 1 0 0 IRF150

.lib nom.lib
.dc lin Vds 0 10 1V Vgs 0 4 0.5V
.probe
.end
